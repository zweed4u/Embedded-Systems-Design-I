filter_mult_inst : filter_mult PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
