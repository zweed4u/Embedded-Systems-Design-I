wave_ram_cos_inst : wave_ram_cos PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
